`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////


module c432_tb;

reg N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
      N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,
      N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,
      N99,N102,N105,N108,N112,N115;
reg [2:0]score;
wire N223,N329,N370,N421,N430,N431,N432;

c432 uut(.N1(N1),.N4(N4),.N11(N11),.N14(N14),.N17(N17),.N21(N21),.N24(N24),.N27(N27),.N30(N30),.N34(N34),.N37(N37),.N40(N40),.N43(N43),.N47(N47),.N50(N50),.N53(N53),.N56(N56),.N60(N60),.N63(N63),.N66(N66),.N69(N69),.N73(N73),.N76(N76),.N79(N79),.N82(N82),.N86(N86),.N89(N89),.N92(N92),.N95(N95),.N99(N99),.N102(N102),.N105(N105),.N108(N108),.N112(N112),.N115(N115),.N223(N223),.N329(N329),.N370(N370),.N421(N421),.N430(N430),.N431(N431),.N432(N432));


initial begin


score <= 3'b000;

//111110000011111000001111100000111110//
N1 <= 1 ; N4 <= 1;  N8 <= 1 ; N11 <= 1 ; N14 <= 1 ; N17 <= 0 ; N21 <= 0;  N24 <= 0 ; N27 <= 0 ; N30 <= 0 ; N34 <= 1 ; N37 <= 1 ;  N40 <=  1; N43 <= 1 ; N47 <= 1 ; N50 <= 0 ; N53 <= 0;  N56 <= 0 ; N60 <= 0 ; N63 <= 0 ; N66 <= 1 ; N69 <= 1;  N73 <= 1 ; N76 <= 1 ; N79 <= 1 ; N82 <= 0 ; N86 <= 0 ; N89 <= 0 ; N92 <= 0 ; N95 <= 0 ; N99 <= 1 ; N102 <= 1 ; N105 <= 1 ; N108 <= 1 ; N112 <= 1 ; N115 <= 0 ;
#10
$display(" input pattern = ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115, "--> golden value = 1001011 "); 
$display(" your answer = " , N223,N329,N370,N421,N430,N431,N432); 
if (N223 == 1'b1 && N329 == 1'b0 && N370 == 1'b0 && N421 == 1'b1 && N430 == 1'b0&& N431 == 1'b1 && N432 == 1'b1 )
begin
	score = score + 3'b001;
end

//110011111111111111110000000000001100//
N1 <= 1 ; N4 <= 1;  N8 <= 0 ; N11 <= 0 ; N14 <= 1 ; N17 <= 1 ; N21 <= 1;  N24 <= 1 ; N27 <= 1 ; N30 <= 1 ; N34 <= 1 ; N37 <= 1 ;  N40 <=  1; N43 <= 1 ; N47 <= 1 ; N50 <= 1 ; N53 <= 1;  N56 <= 1 ; N60 <= 1 ; N63 <= 1 ; N66 <=  0; N69 <= 0;  N73 <= 0 ; N76 <= 0; N79 <= 0 ; N82 <= 0 ; N86 <= 0 ; N89 <= 0 ; N92 <= 0 ; N95 <= 0 ; N99 <= 0 ; N102 <= 0 ; N105 <= 1 ; N108 <= 1 ; N112 <= 0 ; N115 <= 0 ;
#10
$display(" input pattern = ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115," --> golden value = 1111000 "); 
$display(" your answer = ", N223,N329,N370,N421,N430,N431,N432); 
if (N223 == 1'b1 && N329 == 1'b1 && N370 == 1'b1 && N421 == 1'b1 && N430 == 1'b0&& N431 == 1'b0 && N432 == 1'b0 )
begin
	score = score + 3'b001;
end

//000001111111111111110000000000000000//
N1 <= 0 ; N4 <= 0;  N8 <= 0 ; N11 <= 0 ; N14 <= 0 ; N17 <= 1 ; N21 <= 1;  N24 <= 1 ; N27 <= 1 ; N30 <= 1 ; N34 <= 1 ; N37 <= 1 ;  N40 <=  1; N43 <= 1 ; N47 <= 1 ; N50 <= 1 ; N53 <= 1;  N56 <= 1 ; N60 <= 1 ; N63 <= 1 ; N66 <=  0; N69 <= 0;  N73 <= 0 ; N76 <= 0; N79 <= 0 ; N82 <= 0 ; N86 <= 0 ; N89 <= 0 ; N92 <= 0 ; N95 <= 0 ; N99 <= 0 ; N102 <= 0 ; N105 <= 0 ; N108 <= 0 ; N112 <= 0 ; N115 <= 0 ;
#10
$display(" input pattern = ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115," --> golden value = 1001111 "); 
$display(" your answer = ", N223,N329,N370,N421,N430,N431,N432); 
if (N223 == 1'b1 && N329 == 1'b0 && N370 == 1'b0 && N421 == 1'b1 && N430 == 1'b1&& N431 == 1'b1 && N432 == 1'b1 )
begin
	score = score + 3'b001;
end

//000001111111111111110000000000011111//
N1 <= 0 ; N4 <= 0;  N8 <= 0 ; N11 <= 0 ; N14 <= 0 ; N17 <= 1 ; N21 <= 1;  N24 <= 1 ; N27 <= 1 ; N30 <= 1 ; N34 <= 1 ; N37 <= 1 ;  N40 <=  1; N43 <= 1 ; N47 <= 1 ; N50 <= 1 ; N53 <= 1;  N56 <= 1 ; N60 <= 1 ; N63 <= 1 ; N66 <=  0; N69 <= 0;  N73 <= 0 ; N76 <= 0; N79 <= 0 ; N82 <= 0 ; N86 <= 0 ; N89 <= 0 ; N92 <= 0 ; N95 <= 0 ; N99 <= 0 ; N102 <= 1 ; N105 <= 1 ; N108 <= 1 ; N112 <= 1 ; N115 <= 1 ;
#10
$display(" input pattern = ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115," --> golden value = 1001111 "); 
$display(" your answer = ", N223,N329,N370,N421,N430,N431,N432); 
if (N223 == 1'b1 && N329 == 1'b0 && N370 == 1'b0 && N421 == 1'b1 && N430 == 1'b1&& N431 == 1'b1 && N432 == 1'b1 )
begin
	score = score + 3'b001;
end

//111111111111111111001100000000000000//
N1 <= 1 ; N4 <= 1;  N8 <= 1 ; N11 <= 1 ; N14 <= 1 ; N17 <= 1 ; N21 <= 1;  N24 <= 1 ; N27 <= 1 ; N30 <= 1 ; N34 <= 1 ; N37 <= 1 ;  N40 <=  1; N43 <= 1 ; N47 <= 1 ; N50 <= 1 ; N53 <= 1;  N56 <= 1 ; N60 <= 0 ; N63 <= 0 ; N66 <=  1; N69 <= 1;  N73 <= 0 ; N76 <= 0; N79 <= 0 ; N82 <= 0 ; N86 <= 0 ; N89 <= 0 ; N92 <= 0 ; N95 <= 0 ; N99 <= 0 ; N102 <= 0 ; N105 <= 0 ; N108 <= 0 ; N112 <= 0 ; N115 <= 0 ;
#10
$display(" input pattern = ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,N34,N37,N40,N43,N47,N50,N53,N56,N60,N63,N66,N69,N73,N76,N79,N82,N86,N89,N92,N95,N99,N102,N105,N108,N112,N115," --> golden value = 1111011 "); 
$display(" your answer = ", N223,N329,N370,N421,N430,N431,N432); 
if (N223 == 1'b1 && N329 == 1'b1 && N370 == 1'b1 && N421 == 1'b1 && N430 == 1'b0&& N431 == 1'b1 && N432 == 1'b1 )
begin
	score = score + 3'b001;
end

if (score == 3'b101)
begin
$display("You're all correct!!!");
$display("  ***    *** ");
$display(" *****  *****");
$display("**************");
$display(" ************ ");
$display("  **********  ");
$display("   ********   ");
$display("    ******    ");
$display("     ****     ");
$display("      **      ");
end
else
$display("WRONG");
end
  
endmodule