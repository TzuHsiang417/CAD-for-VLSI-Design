`timescale 1ns / 1ps


module c880_tb;

reg N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,
      N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,
      N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,
      N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,
      N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,
      N219,N228,N237,N246,N255,N259,N260,N261,N267,N268;
	  
reg [2:0]score;
wire N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,
       N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,
       N865,N866,N874,N878,N879,N880;

c880 uut(.N1(N1),.N8(N8),.N13(N13),.N17(N17),.N26(N26),.N29(N29),.N36(N36),.N42(N42),.N51(N51),.N55(N55),.
      N59(N59),.N68(N68),.N72(N72),.N73(N73),.N74(N74),.N75(N75),.N80(N80),.N85(N85),.N86(N86),.N87(N87),.
      N88(N88),.N89(N89),.N90(N90),.N91(N91),.N96(N96),.N101(N101),.N106(N106),.N111(N111),.N116(N116),.N121(N121),.
      N126(N126),.N130(N130),.N135(N135),.N138(N138),.N143(N143),.N146(N146),.N149(N149),.N152(N152),.N153(N153),.N156(N156),.
      N159(N159),.N165(N165),.N171(N171),.N177(N177),.N183(N183),.N189(N189),.N195(N195),.N201(N201),.N207(N207),.N210(N210),.
      N219(N219),.N228(N228),.N237(N237),.N246(N246),.N255(N255),.N259(N259),.N260(N260),.N261(N261),.N267(N267),.N268(N268),.N388(N388),.N389(N389),.N390(N390),.N391(N391),.N418(N418),.N419(N419),.N420(N420),.N421(N421),.N422(N422),.N423(N423),.
      N446(N446),.N447(N447),.N448(N448),.N449(N449),.N450(N450),.N767(N767),.N768(N768),.N850(N850),.N863(N863),.N864(N864),.
      N865(N865),.N866(N866),.N874(N874),.N878(N878),.N879(N879),.N880(N880));




initial begin


score <= 3'b000;

//001100011111001110000000001111111111111111100001111111111000//
N1 <= 0 ; N8 <= 0 ; N13 <= 1 ; N17 <= 1 ; N26 <= 0 ; N29 <= 0 ; N36 <= 0 ; N42 <= 1 ; N51 <= 1 ; N55 <= 1 ; N59 <= 1 ; N68 <= 1 ; N72 <= 0 ; N73 <= 0 ; N74 <= 1 ; N75 <= 1 ; N80 <= 1 ; N85 <= 0 ; N86 <= 0 ; N87 <= 0 ; N88 <= 0 ; N89 <= 0 ; N90 <= 0 ; N91 <= 0 ; N96 <= 0 ; N101 <= 0 ; N106 <= 1 ; N111 <= 1 ; N116 <= 1 ; N121 <= 1 ; N126 <= 1 ; N130 <= 1 ; N135 <= 1 ; N138 <= 1 ; N143 <= 1 ; N146 <= 1 ; N149 <= 1 ; N152 <= 1 ; N153 <= 1 ; N156 <= 1 ; N159 <= 1 ; N165 <= 1 ; N171 <= 1 ; N177 <= 0 ; N183 <= 0 ; N189 <= 0 ; N195 <= 0 ; N201 <= 1 ; N207 <= 1 ; N210 <= 1 ; N219 <= 1 ; N228 <= 1 ; N237 <= 1 ; N246 <= 1 ; N255 <= 1 ; N259 <= 1 ; N260 <= 1 ; N261 <= 0 ; N267 <= 0 ; N268 <= 0;
#10
$display(" input pattern = " ,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268," --> golden value = 00000101101000010111111111"); 
$display(" your answer = " ,N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880); 
if (N388 == 1'b0 && N389 == 1'b0 && N390 == 1'b0 && N391 == 1'b0 && N418 == 1'b0 && N419 == 1'b1 && N420 == 1'b0 && N421 == 1'b1 && N422 == 1'b1 && N423 == 1'b0 && N446 == 1'b1 && N447 == 1'b0 && N448 == 1'b0 && N449 == 1'b0 && N450 == 1'b0 && N767 == 1'b1 && N768 == 1'b0 && N850 == 1'b1 && N863 == 1'b1 && N864 == 1'b1 && N865 == 1'b1 && N866 == 1'b1 && N874 == 1'b1 && N878 == 1'b1 && N879 == 1'b1 && N880 == 1'b1 )
begin
	score = score + 3'b001;
end

//111000000001110001111111111111111110000000111111111110001111//
N1 <= 1 ; N8 <= 1 ; N13 <= 1 ; N17 <= 0 ; N26 <= 0 ; N29 <= 0 ; N36 <= 0 ; N42 <= 0 ; N51 <= 0 ; N55 <= 0 ; N59 <= 0 ; N68 <= 1 ; N72 <= 1 ; N73 <= 1 ; N74 <= 0 ; N75 <= 0 ; N80 <= 0 ; N85 <= 1 ; N86 <= 1 ; N87 <= 1 ; N88 <= 1 ; N89 <= 1 ; N90 <= 1 ; N91 <= 1 ; N96 <= 1 ; N101 <= 1 ; N106 <= 1 ; N111 <= 1 ; N116 <= 1 ; N121 <= 1 ; N126 <= 1 ; N130 <= 1 ; N135 <= 1 ; N138 <= 1 ; N143 <= 1 ; N146 <= 0 ; N149 <= 0 ; N152 <= 0 ; N153 <= 0 ; N156 <= 0 ; N159 <= 0 ; N165 <= 0 ; N171 <= 1 ; N177 <= 1 ; N183 <= 1 ; N189 <= 1 ; N195 <= 1 ; N201 <= 1 ; N207 <= 1 ; N210 <= 1 ; N219 <= 1 ; N228 <= 1 ; N237 <= 1 ; N246 <= 0 ; N255 <= 0 ; N259 <= 0 ; N260 <= 1 ; N261 <= 1 ; N267 <= 1 ; N268 <= 1;
#10
$display(" input pattern = " ,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268," --> golden value = 00010111111000100111101111"); 
$display(" your answer = ", N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880); 
if (N388 == 1'b0 && N389 == 1'b0 && N390 == 1'b0 && N391 == 1'b1 && N418 == 1'b0 && N419 == 1'b1 && N420 == 1'b1 && N421 == 1'b1 && N422 == 1'b1 && N423 == 1'b1 && N446 == 1'b1 && N447 == 1'b0 && N448 == 1'b0 && N449 == 1'b0 && N450 == 1'b1 && N767 == 1'b0 && N768 == 1'b0 && N850 == 1'b1 && N863 == 1'b1 && N864 == 1'b1 && N865 == 1'b1 && N866 == 1'b0 && N874 == 1'b1 && N878 == 1'b1 && N879 == 1'b1 && N880 == 1'b1 )
begin
	score = score + 3'b001;
end
 
//000011111111111111111000000000000000011111111111111110000011//
N1 <= 0 ; N8 <= 0 ; N13 <= 0 ; N17 <= 0 ; N26 <= 1 ; N29 <= 1 ; N36 <= 1 ; N42 <= 1 ; N51 <= 1 ; N55 <= 1 ; N59 <= 1 ; N68 <= 1 ; N72 <= 1 ; N73 <= 1 ; N74 <= 1 ; N75 <= 1 ; N80 <= 1 ; N85 <= 1 ; N86 <= 1 ; N87 <= 1 ; N88 <= 1 ; N89 <= 0 ; N90 <= 0 ; N91 <= 0 ; N96 <= 0 ; N101 <= 0 ; N106 <= 0 ; N111 <= 0 ; N116 <= 0 ; N121 <= 0 ; N126 <= 0 ; N130 <= 0 ; N135 <= 0 ; N138 <= 0 ; N143 <= 0 ; N146 <= 0 ; N149 <= 0 ; N152 <= 1 ; N153 <= 1 ; N156 <= 1 ; N159 <= 1 ; N165 <= 1 ; N171 <= 1 ; N177 <= 1 ; N183 <= 1 ; N189 <= 1 ; N195 <= 1 ; N201 <= 1 ; N207 <= 1 ; N210 <= 1 ; N219 <= 1 ; N228 <= 1 ; N237 <= 1 ; N246 <= 0 ; N255 <= 0 ; N259 <= 0 ; N260 <= 0 ; N261 <= 0 ; N267 <= 1 ; N268 <= 1;
#10
$display(" input pattern = " ,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268," --> golden value = 11110100001000001111111111"); 
$display(" your answer = ", N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880); 
if (N388 == 1'b1 && N389 == 1'b1 && N390 == 1'b1 && N391 == 1'b1 && N418 == 1'b0 && N419 == 1'b1 && N420 == 1'b0 && N421 == 1'b0 && N422 == 1'b0 && N423 == 1'b0 && N446 == 1'b1 && N447 == 1'b0 && N448 == 1'b0 && N449 == 1'b0 && N450 == 1'b0 && N767 == 1'b0 && N768 == 1'b1 && N850 == 1'b1 && N863 == 1'b1 && N864 == 1'b1 && N865 == 1'b1 && N866 == 1'b1 && N874 == 1'b1 && N878 == 1'b1 && N879 == 1'b1 && N880 == 1'b1 )
begin
	score = score + 3'b001;
end

//000000000000000000000000000000000000000000000000000000000000//
N1 <= 0 ; N8 <= 0 ; N13 <= 0 ; N17 <= 0 ; N26 <= 0 ; N29 <= 0 ; N36 <= 0 ; N42 <= 0 ; N51 <= 0 ; N55 <= 0 ; N59 <= 0 ; N68 <= 0 ; N72 <= 0 ; N73 <= 0 ; N74 <= 0 ; N75 <= 0 ; N80 <= 0 ; N85 <= 0 ; N86 <= 0 ; N87 <= 0 ; N88 <= 0 ; N89 <= 0 ; N90 <= 0 ; N91 <= 0 ; N96 <= 0 ; N101 <= 0 ; N106 <= 0 ; N111 <= 0 ; N116 <= 0 ; N121 <= 0 ; N126 <= 0 ; N130 <= 0 ; N135 <= 0 ; N138 <= 0 ; N143 <= 0 ; N146 <= 0 ; N149 <= 0 ; N152 <= 0 ; N153 <= 0 ; N156 <= 0 ; N159 <= 0 ; N165 <= 0 ; N171 <= 0 ; N177 <= 0 ; N183 <= 0 ; N189 <= 0 ; N195 <= 0 ; N201 <= 0 ; N207 <= 0 ; N210 <= 0 ; N219 <= 0 ; N228 <= 0 ; N237 <= 0 ; N246 <= 0 ; N255 <= 0 ; N259 <= 0 ; N260 <= 0 ; N261 <= 0 ; N267 <= 0 ; N268 <= 0;
#10
$display(" input pattern = " ,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268," --> golden value = 00000111101000000000000000"); 
$display(" your answer = ", N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880); 
if (N388 == 1'b0 && N389 == 1'b0 && N390 == 1'b0 && N391 == 1'b0 && N418 == 1'b0 && N419 == 1'b1 && N420 == 1'b1 && N421 == 1'b1 && N422 == 1'b1 && N423 == 1'b0 && N446 == 1'b1 && N447 == 1'b0 && N448 == 1'b0 && N449 == 1'b0 && N450 == 1'b0 && N767 == 1'b0 && N768 == 1'b0 && N850 == 1'b0 && N863 == 1'b0 && N864 == 1'b0 && N865 == 1'b0 && N866 == 1'b0 && N874 == 1'b0 && N878 == 1'b0 && N879 == 1'b0 && N880 == 1'b0 )
begin
	score = score + 3'b001;
end

//111111111111111111111111111111111111111111111111111111111111//
N1 <= 1 ; N8 <= 1 ; N13 <= 1 ; N17 <= 1 ; N26 <= 1 ; N29 <= 1 ; N36 <= 1 ; N42 <= 1 ; N51 <= 1 ; N55 <= 1 ; N59 <= 1 ; N68 <= 1 ; N72 <= 1 ; N73 <= 1 ; N74 <= 1 ; N75 <= 1 ; N80 <= 1 ; N85 <= 1 ; N86 <= 1 ; N87 <= 1 ; N88 <= 1 ; N89 <= 1 ; N90 <= 1 ; N91 <= 1 ; N96 <= 1 ; N101 <= 1 ; N106 <= 1 ; N111 <= 1 ; N116 <= 1 ; N121 <= 1 ; N126 <= 1 ; N130 <= 1 ; N135 <= 1 ; N138 <= 1 ; N143 <= 1 ; N146 <= 1 ; N149 <= 1 ; N152 <= 1 ; N153 <= 1 ; N156 <= 1 ; N159 <= 1 ; N165 <= 1 ; N171 <= 1 ; N177 <= 1 ; N183 <= 1 ; N189 <= 1 ; N195 <= 1 ; N201 <= 1 ; N207 <= 1 ; N210 <= 1 ; N219 <= 1 ; N228 <= 1 ; N237 <= 1 ; N246 <= 1 ; N255 <= 1 ; N259 <= 1 ; N260 <= 1 ; N261 <= 1 ; N267 <= 1 ; N268 <= 1;
#10
$display(" input pattern = " ,N1,N8,N13,N17,N26,N29,N36,N42,N51,N55,N59,N68,N72,N73,N74,N75,N80,N85,N86,N87,N88,N89,N90,N91,N96,N101,N106,N111,N116,N121,N126,N130,N135,N138,N143,N146,N149,N152,N153,N156,N159,N165,N171,N177,N183,N189,N195,N201,N207,N210,N219,N228,N237,N246,N255,N259,N260,N261,N267,N268," --> golden value = 11111100010111100111111111"); 
$display(" your answer = ", N388,N389,N390,N391,N418,N419,N420,N421,N422,N423,N446,N447,N448,N449,N450,N767,N768,N850,N863,N864,N865,N866,N874,N878,N879,N880); 
if (N388 == 1'b1 && N389 == 1'b1 && N390 == 1'b1 && N391 == 1'b1 && N418 == 1'b1 && N419 == 1'b1 && N420 == 1'b0 && N421 == 1'b0 && N422 == 1'b0 && N423 == 1'b1 && N446 == 1'b0 && N447 == 1'b1 && N448 == 1'b1 && N449 == 1'b1 && N450 == 1'b1 && N767 == 1'b0 && N768 == 1'b0 && N850 == 1'b1 && N863 == 1'b1 && N864 == 1'b1 && N865 == 1'b1 && N866 == 1'b1 && N874 == 1'b1 && N878 == 1'b1 && N879 == 1'b1 && N880 == 1'b1 )
begin
	score = score + 3'b001;
end

if (score == 3'b101)
begin
$display("You're all correct!!!");
$display("  ***    *** ");
$display(" *****  *****");
$display("**************");
$display(" ************ ");
$display("  **********  ");
$display("   ********   ");
$display("    ******    ");
$display("     ****     ");
$display("      **      ");
end
else
$display("WRONG");
end
  
endmodule